
no_st_flush: assume property(##2 core.id_unit.st_flush_i == 0);
